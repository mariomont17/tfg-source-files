`ifndef BUS_ENV_PKG_SV
`define BUS_ENV_PKG_SV
`include "uvm_macros.svh"
package bus_env_pkg;
  import uvm_pkg::*;
	`include "bus_seq_item.sv"
	`include "bus_sqr.sv"
	`include "bus_driver.sv"
	`include "bus_monitor.sv"
	`include "bus_agent.sv"
	`include "bus_scoreboard.sv"
	`include "bus_coverage.sv"
	`include "bus_env.sv"
endpackage : bus_env_pkg
`endif
