`include "uvm_macros.svh"
package bus_top_pkg;
	`include "bus_interface.sv"
	`include "bus_env_pkg.sv"
	`include "bus_seq_pkg.sv"
	`include "bus_test_pkg.sv"
endpackage : bus_top_pkg
